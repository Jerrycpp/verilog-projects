module debounce (clk, inp, out, rst);
    input clk, inp, rst;
    output out;
endmodule