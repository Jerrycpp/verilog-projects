module slave_i2c_tb;
    reg clk;

    wire sda, scl;
    

endmodule